magic
tech scmos
magscale 1 2
timestamp 1498914250
<< metal1 >>
rect 493 143 499 156
rect 413 137 435 143
rect 477 137 499 143
rect 532 137 547 143
rect 509 117 531 123
<< m2contact >>
rect 188 156 196 164
rect 492 156 500 164
rect 556 156 564 164
rect 12 136 20 144
rect 348 136 356 144
rect 364 138 372 146
rect 524 136 532 144
rect 44 116 52 124
rect 188 118 196 126
rect 268 116 276 124
rect 316 116 324 124
rect 332 116 340 124
rect 364 116 372 124
rect 396 116 404 124
rect 460 116 468 124
rect 284 96 292 104
rect 60 76 68 84
rect 436 76 444 84
<< metal2 >>
rect 189 237 211 243
rect 189 164 195 237
rect 13 124 19 136
rect 189 126 195 136
rect 269 124 275 243
rect 317 124 323 243
rect 189 117 195 118
rect 45 103 51 116
rect 45 97 67 103
rect 61 84 67 97
rect 349 84 355 136
rect 397 124 403 136
rect 461 124 467 243
rect 493 237 515 243
rect 493 164 499 237
rect 493 124 499 156
rect 365 104 371 116
rect 445 -23 451 76
<< m3contact >>
rect 188 136 196 144
rect 12 116 20 124
rect 364 138 372 144
rect 364 136 372 138
rect 396 136 404 144
rect 332 116 340 124
rect 284 96 292 104
rect 556 156 564 164
rect 524 136 532 144
rect 492 116 500 124
rect 364 96 372 104
rect 348 76 356 84
rect 444 76 452 84
<< metal3 >>
rect 564 157 595 163
rect 196 137 364 143
rect 404 137 524 143
rect -19 117 12 123
rect 340 117 492 123
rect 292 97 364 103
rect 356 77 444 83
use BUFX2  BUFX2_1
timestamp 1498914250
transform -1 0 56 0 -1 210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_1
timestamp 1498914250
transform -1 0 248 0 -1 210
box 0 0 192 200
use MUX2X1  MUX2X1_1
timestamp 1498914250
transform -1 0 344 0 -1 210
box 0 0 96 200
use OAI22X1  OAI22X1_1
timestamp 1498914250
transform -1 0 424 0 -1 210
box 0 0 80 200
use OAI21X1  OAI21X1_1
timestamp 1498914250
transform -1 0 488 0 -1 210
box 0 0 64 200
use INVX1  INVX1_1
timestamp 1498914250
transform 1 0 488 0 -1 210
box 0 0 32 200
use NOR2X1  NOR2X1_1
timestamp 1498914250
transform -1 0 568 0 -1 210
box 0 0 48 200
<< labels >>
flabel metal3 592 160 592 160 3 FreeSans 24 0 0 0 i1
flabel metal2 464 240 464 240 3 FreeSans 24 90 0 0 i2
flabel metal2 272 240 272 240 3 FreeSans 24 90 0 0 i3
flabel metal2 320 240 320 240 3 FreeSans 24 90 0 0 i4
flabel metal2 448 -20 448 -20 7 FreeSans 24 270 0 0 sel<0>
flabel metal2 512 240 512 240 3 FreeSans 24 90 0 0 sel<1>
flabel metal2 208 240 208 240 3 FreeSans 24 90 0 0 clk
flabel metal3 -16 120 -16 120 7 FreeSans 24 0 0 0 out
<< end >>
